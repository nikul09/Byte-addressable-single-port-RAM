
`ifndef ram_define_sv
`define ram_define_sv

`define addr_width 5
`define data_width 32
`define mem_depth 32

`endif
