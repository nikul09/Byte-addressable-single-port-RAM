
`include "define.sv" 

package ram_pkg;


`include "transection.sv"
`include "my_config_db.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "schoreboard.sv"
`include "agent.sv"
`include "environment.sv"
`include "test.sv"

endpackage
